`default_nettype 

module segment_logic (
    input wire clk,
    input wire rst_n,
    input wire 
);
    
endmodule